----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 07/22/2024 12:07:06 PM
-- Design Name: 
-- Module Name: tanh_lut - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity tanh_lut is
    Port (
        clka    : in  STD_LOGIC;
        ena     : in  STD_LOGIC;
        addra   : in  STD_LOGIC_VECTOR (7 downto 0);
        douta   : out STD_LOGIC_VECTOR (31 downto 0)
    );
end tanh_lut;

architecture Behavioral of tanh_lut is

    type memory_array is array (0 to 255) of STD_LOGIC_VECTOR(31 downto 0);
    constant tanh_lut : memory_array := (
        X"00000000",
        X"0003FFEA",
        X"0007FF55",
        X"000BFDC0",
        X"000FFAAC",
        X"0013F59B",
        X"0017EE10",
        X"001BE38D",
        X"001FD599",
        X"0023C3BA",
        X"0027AD78",
        X"002B9260",
        X"002F71FF",
        X"00334BE3",
        X"00371FA0",
        X"003AECCB",
        X"003EB2FD",
        X"004271D1",
        X"004628E6",
        X"0049D7DF",
        X"004D7E62",
        X"00511C19",
        X"0054B0B1",
        X"00583BDC",
        X"005BBD4F",
        X"005F34C4",
        X"0062A1F8",
        X"006604AC",
        X"00695CA7",
        X"006CA9B2",
        X"006FEB9A",
        X"00732232",
        X"00764D4F",
        X"00796CCB",
        X"007C8084",
        X"007F885B",
        X"00828437",
        X"00857400",
        X"008857A3",
        X"008B2F12",
        X"008DFA3F",
        X"0090B922",
        X"00936BB7",
        X"009611FB",
        X"0098ABEF",
        X"009B3998",
        X"009DBAFC",
        X"00A03025",
        X"00A2991F",
        X"00A4F5F9",
        X"00A746C4",
        X"00A98B94",
        X"00ABC47F",
        X"00ADF19C",
        X"00B01304",
        X"00B228D4",
        X"00B43328",
        X"00B6321F",
        X"00B825D8",
        X"00BA0E77",
        X"00BBEC1C",
        X"00BDBEEC",
        X"00BF870D",
        X"00C144A3",
        X"00C2F7D5",
        X"00C4A0CB",
        X"00C63FAE",
        X"00C7D4A5",
        X"00C95FD9",
        X"00CAE175",
        X"00CC59A3",
        X"00CDC88C",
        X"00CF2E5A",
        X"00D08B3A",
        X"00D1DF54",
        X"00D32AD5",
        X"00D46DE5",
        X"00D5A8B1",
        X"00D6DB62",
        X"00D80623",
        X"00D9291D",
        X"00DA447B",
        X"00DB5865",
        X"00DC6506",
        X"00DD6A85",
        X"00DE690A",
        X"00DF60BF",
        X"00E051CA",
        X"00E13C52",
        X"00E2207E",
        X"00E2FE74",
        X"00E3D658",
        X"00E4A851",
        X"00E57482",
        X"00E63B10",
        X"00E6FC1C",
        X"00E7B7CB",
        X"00E86E3E",
        X"00E91F96",
        X"00E9CBF5",
        X"00EA737A",
        X"00EB1645",
        X"00EBB475",
        X"00EC4E28",
        X"00ECE37D",
        X"00ED7490",
        X"00EE017E",
        X"00EE8A63",
        X"00EF0F5A",
        X"00EF907F",
        X"00F00DEA",
        X"00F087B6",
        X"00F0FDFC",
        X"00F170D5",
        X"00F1E057",
        X"00F24C9B",
        X"00F2B5B7",
        X"00F31BC2",
        X"00F37ED1",
        X"00F3DEF9",
        X"00F43C4F",
        X"00F496E7",
        X"00F4EED5",
        X"00F5442C",
        X"00F596FF",
        X"00F5E75F",
        X"00F6355F",
        X"00F68110",
        X"00F6CA82",
        X"00F711C7",
        X"00F756ED",
        X"00F79A05",
        X"00F7DB1E",
        X"00F81A45",
        X"00F8578B",
        X"00F892FC",
        X"00F8CCA6",
        X"00F90497",
        X"00F93ADB",
        X"00F96F7F",
        X"00F9A28F",
        X"00F9D416",
        X"00FA0420",
        X"00FA32B9",
        X"00FA5FEB",
        X"00FA8BC1",
        X"00FAB644",
        X"00FADF80",
        X"00FB077D",
        X"00FB2E45",
        X"00FB53E2",
        X"00FB785C",
        X"00FB9BBB",
        X"00FBBE08",
        X"00FBDF4C",
        X"00FBFF8E",
        X"00FC1ED5",
        X"00FC3D2A",
        X"00FC5A94",
        X"00FC7719",
        X"00FC92C1",
        X"00FCAD91",
        X"00FCC791",
        X"00FCE0C7",
        X"00FCF939",
        X"00FD10EC",
        X"00FD27E7",
        X"00FD3E2F",
        X"00FD53C9",
        X"00FD68BB",
        X"00FD7D09",
        X"00FD90B9",
        X"00FDA3D0",
        X"00FDB651",
        X"00FDC842",
        X"00FDD9A7",
        X"00FDEA84",
        X"00FDFADE",
        X"00FE0AB7",
        X"00FE1A15",
        X"00FE28FA",
        X"00FE376B",
        X"00FE456B",
        X"00FE52FE",
        X"00FE6026",
        X"00FE6CE7",
        X"00FE7945",
        X"00FE8541",
        X"00FE90E0",
        X"00FE9C24",
        X"00FEA70F",
        X"00FEB1A5",
        X"00FEBBE8",
        X"00FEC5DB",
        X"00FECF7F",
        X"00FED8D8",
        X"00FEE1E8",
        X"00FEEAB0",
        X"00FEF334",
        X"00FEFB75",
        X"00FF0375",
        X"00FF0B36",
        X"00FF12BB",
        X"00FF1A04",
        X"00FF2115",
        X"00FF27EE",
        X"00FF2E91",
        X"00FF3500",
        X"00FF3B3C",
        X"00FF4148",
        X"00FF4724",
        X"00FF4CD2",
        X"00FF5253",
        X"00FF57A9",
        X"00FF5CD5",
        X"00FF61D9",
        X"00FF66B5",
        X"00FF6B6B",
        X"00FF6FFC",
        X"00FF7469",
        X"00FF78B4",
        X"00FF7CDC",
        X"00FF80E4",
        X"00FF84CC",
        X"00FF8896",
        X"00FF8C41",
        X"00FF8FD0",
        X"00FF9343",
        X"00FF969B",
        X"00FF99D8",
        X"00FF9CFC",
        X"00FFA008",
        X"00FFA2FB",
        X"00FFA5D7",
        X"00FFA89D",
        X"00FFAB4D",
        X"00FFADE7",
        X"00FFB06D",
        X"00FFB2E0",
        X"00FFB53F",
        X"00FFB78B",
        X"00FFB9C6",
        X"00FFBBEF",
        X"00FFBE06",
        X"00FFC00E",
        X"00FFC205",
        X"00FFC3ED",
        X"00FFC5C6",
        X"00FFC790",
        X"00FFC94D",
        X"00FFCAFB",
        X"00FFCC9D",
        X"00FFCE31",
        X"00FFCFB9",
        X"00FFD136",
        X"00FFD2A6"
    );

    signal addr_reg1, addr_reg2 : STD_LOGIC_VECTOR(7 downto 0);
    signal data_reg1, data_reg2 : STD_LOGIC_VECTOR(31 downto 0);

begin
    process(clka)
    begin
        if rising_edge(clka) then
            if ena = '1' then
                addr_reg1 <= addra;
                data_reg1 <= tanh_lut(to_integer(unsigned(addra)));
                addr_reg2 <= addr_reg1;
                data_reg2 <= data_reg1;
            end if;
        end if;
    end process;

    douta <= data_reg2;

end Behavioral;